`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: MIT
// Engineer: Schuyler Senft-Grupp
// 
// Create Date:    14:30:37 07/04/2014 
// Design Name: 
// Module Name:    DataStorageAcc 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module DataStorageAcc(
    input [31:0] DataIn,
    output reg [7:0] DataOut,
    input FastTrigger,
    input ReadEnable,
    input WriteClock,
    input ReadClock,
    input Reset,
    output reg DataReady = 0,
	 output [7:0] gDataOut,
	 output reg GenStrobe = 0
    );


	reg byteNumber; //read high (1) or low byte (0) 
	reg [3:0] fifoNumber = 4'b0001;
	reg [7:0] GenDataOut = 8'b0;
	wire [15:0] dataOutDQD;
	wire [15:0] dataOutDID;
	wire [15:0] dataOutDQ;
	wire [15:0] dataOutDI;
	
	reg [10:0] readCounts = 11'd0; //this is 10 bits - 512 data points * 2 bytes each
	
	assign gDataOut = GenDataOut;
	
	
	wire sendEOD = (readCounts == 11'd1024);
	//state machine for sending "end-of-data" bytes
	parameter WAIT_FOR_END  = 4'b0001;
	parameter END1				= 4'b0010;
	parameter PAUSE 			= 4'b0100;
	parameter END2				= 4'b1000;
	
	//TO DO I should probably implement 4 end bytes with the 3rd and 4th the opposite order of 1 and 2
	
	(* FSM_ENCODING="ONE-HOT", SAFE_IMPLEMENTATION="NO" *) reg [3:0] eofState = WAIT_FOR_END;
	always@(posedge ReadClock) begin
		(* FULL_CASE, PARALLEL_CASE *) case (eofState)
		WAIT_FOR_END:begin
			GenStrobe <= 1'b0;
			GenDataOut <= 8'b00000000;
			if(sendEOD)
				eofState <= END1;
			else
				eofState <= WAIT_FOR_END;
		end
		END1: begin
			eofState <= PAUSE;
			GenDataOut <= 8'b10000000;
			GenStrobe <= 1'b1;
		end
		PAUSE:begin
			eofState <= END2;
			GenDataOut <= 8'b00000000;
			GenStrobe <= 1'b0;
		end
		END2: begin
			eofState <= WAIT_FOR_END;
			GenDataOut <= 8'b00000001;
			GenStrobe <= 1'b1;
		end
		endcase
	end
	
	
	parameter WAIT_TO_TRANSMIT = 5'b00001;
	parameter DQD_READ		= 5'b00010;
	parameter DID_READ		= 5'b00100;
	parameter DQ_READ			= 5'b01000;
	parameter DI_READ 		= 5'b10000;
	
	
	//Wait until data is available on all fifos
	wire dataReadyFromAcc = dataReadyToReadDI | dataReadyToReadDID | dataReadyToReadDQ | dataReadyToReadDQD;
	
	
	always@(posedge ReadClock) begin
		DataReady <= (state != WAIT_TO_TRANSMIT);
		if(state == WAIT_TO_TRANSMIT) begin
			byteNumber <= 0;
			readCounts <= 0;
		end
		else if (ReadEnable) begin
			byteNumber <= ~byteNumber;
			readCounts <= readCounts + 1;
		end
	end
	
	reg dqRd = 0, dqdRd = 0, diRd = 0, didRd = 0;
	
	wire fsmReset = (readCounts == 11'd1024) | Reset;  //1024
	
	//note: the read signals should only pulse high for 1 clock cycle
	//after the current data has already been read
	
	(* FSM_ENCODING="ONE-HOT", SAFE_IMPLEMENTATION="NO" *) reg [4:0] state = WAIT_TO_TRANSMIT;
	always@(posedge ReadClock)
      if (fsmReset) begin
         state <= WAIT_TO_TRANSMIT;
      end
      else
         (* FULL_CASE, PARALLEL_CASE *) case (state)
			WAIT_TO_TRANSMIT: begin
				dqRd  <= 0;
				dqdRd <= 0;
				diRd  <= 0;
				didRd <= 0;
				if(dataReadyFromAcc)
					state <= DQD_READ;
				else
					state <=WAIT_TO_TRANSMIT;
			end
			DQD_READ: begin
				dqRd  <= 0;
				diRd  <= 0;
				didRd <= 0;
				if(ReadEnable & (byteNumber)) begin
					state <= DID_READ;
					dqdRd <= 1;
				end
				else begin
					state <=DQD_READ;
					dqdRd <= 0;
				end
				if(byteNumber)
					DataOut <= dataOutDQD[7:0];
				else
					DataOut <= dataOutDQD[15:8];				
			end
			DID_READ: begin
				dqdRd <= 0;
				dqRd  <= 0;
				diRd <= 0;
				if(ReadEnable & (byteNumber)) begin
					state <= DQ_READ;
					didRd <= 1;
				end
				else begin
					state <=DID_READ;
					didRd <= 0;
				end
				if(byteNumber)
					DataOut <= dataOutDID[7:0];
				else
					DataOut <= dataOutDID[15:8];				
			end			
			DQ_READ: begin
				dqdRd <= 0;
				diRd  <= 0;
				didRd <= 0;
				
				if(ReadEnable & (byteNumber)) begin
					state <= DI_READ;
					dqRd <= 1;
				end
				else begin
					state <=DQ_READ;
					dqRd <= 0;
				end
				
				if(byteNumber)
					DataOut <= dataOutDQ[7:0];
				else
					DataOut <= dataOutDQ[15:8];
			end
			DI_READ: begin
				dqdRd <= 0;
				dqRd  <= 0;
				didRd <= 0;
				
				if(ReadEnable & (byteNumber)) begin
					state <= DQD_READ;	//move to next state
					diRd <= 1;
				end
				else begin
					state <=DI_READ; 	//stay at this state
					diRd <= 0;
				end
				
				if(byteNumber)
					DataOut <= dataOutDI[7:0];
				else
					DataOut <= dataOutDI[15:8];
			end
		endcase
			
			
//fifos 
DataAccumulator DI (
    .clk(WriteClock),
    .clkSlow(ReadClock), 
    .inputData(DataIn[31:24]), 
    .dataCaptureStrobe(FastTrigger), 
    .dataRead(diRd), 
    .rst(Reset), 
    .dataReadyToRead(dataReadyToReadDI), 
    .dataEmpty(dataEmptyDI), 
    .dataOut(dataOutDI)
    );
	 
DataAccumulator DID (
    .clk(WriteClock),
    .clkSlow(ReadClock), 
    .inputData(DataIn[23:16]), 
    .dataCaptureStrobe(FastTrigger), 
    .dataRead(didRd), 
    .rst(Reset), 
    .dataReadyToRead(dataReadyToReadDID), 
    .dataEmpty(dataEmptyDID), 
    .dataOut(dataOutDID)
    );
	 
DataAccumulator DQ (
    .clk(WriteClock),
    .clkSlow(ReadClock), 
    .inputData(DataIn[15:8]), 
    .dataCaptureStrobe(FastTrigger), 
    .dataRead(dqRd), 
    .rst(Reset), 
    .dataReadyToRead(dataReadyToReadDQ), 
    .dataEmpty(dataEmptyDQ), 
    .dataOut(dataOutDQ)
    );
	 
DataAccumulator DQD (
    .clk(WriteClock),
    .clkSlow(ReadClock), 
    .inputData(DataIn[7:0]), 
    .dataCaptureStrobe(FastTrigger), 
    .dataRead(dqdRd), 
    .rst(Reset), 
    .dataReadyToRead(dataReadyToReadDQD), 
    .dataEmpty(dataEmptyDQD), 
    .dataOut(dataOutDQD)
    );
	 

endmodule
